*                                               Revised: Monday, October 30, 2017
* E:\ORCAD\SOILDERSTATION\ORCAD_HAKKO.DSN       Revision: 
* 
* 
* 
* 
* 
VCC 15001 0 
U1 14994 14995 14989 15001 0    LM358
U2 14992 14990 14997 14991 14989 15001 0 14993 ATtiny13
U3 15004 15001 0 7805
R1 14995 14989 100K
R2 15001 14988 2K7
U4 15001 14991 0 50K
R3 14988 14994 10K
R4 14995 0 10K
R5 14997 14999 1K
R6 14996 0 10K
R7 14996 15000 10K
R8 15005 15003 1K5
R9 15002 0 390
C1 14988 0 102
C2 15004 0 1000uF
C3 15001 0 100uF
R10 15001 14993 10K
R11 0 16024 1M
J1 15004 0 DC Jack
J2 14988 16024 0 SENSOR
J3 15001 14992 14990 0 DISPLAY
J4 15003 15004 HEATER
D1 15001 15002 GREEN
D2 15004 15005 RED
SW1 0 14993 BUTTON
Q1 14999 15001 14996 A1015
Q2 15003 15000 0 IRF540N/TO
.END
